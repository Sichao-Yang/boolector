// Note: The license below is based on the template at:
// http://opensource.org/licenses/BSD-3-Clause
// Copyright (C) 2020 Regents of the University of Texas
//All rights reserved.

// Redistribution and use in source and binary forms, with or without
// modification, are permitted provided that the following conditions are
// met:

// o Redistributions of source code must retain the above copyright
//   notice, this list of conditions and the following disclaimer.

// o Redistributions in binary form must reproduce the above copyright
//   notice, this list of conditions and the following disclaimer in the
//   documentation and/or other materials provided with the distribution.

// o Neither the name of the copyright holders nor the names of its
//   contributors may be used to endorse or promote products derived
//   from this software without specific prior written permission.

// THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS
// "AS IS" AND ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT
// LIMITED TO, THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR
// A PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT
// HOLDER OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT, INDIRECT, INCIDENTAL,
// SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES (INCLUDING, BUT NOT
// LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES; LOSS OF USE,
// DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER CAUSED AND ON ANY
// THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT
// (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE
// OF THIS SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.

// Original Author(s):
// Mertcan Temel         <mert@utexas.edu>

// DO NOT REMOVE:
// This file is generated by Temel's multiplier generator. Download from https://github.com/temelmertcan/multgen.

// Specification module to help understand what the design implements.
module WT_USP_RP_2x2_noX_spec (
        input logic [1:0] IN1,
        input logic [1:0] IN2,
        input logic [0:0] IN3, //redundant
        output logic design_is_correct, // is set to 1 iff the output of WT_USP_RP_2x2_noX matches its spec.
        output logic [3:0] design_res,
        output logic [3:0] spec_res);
    
    assign spec_res = unsigned'(IN1) * unsigned'(IN2);
    WT_USP_RP_2x2_noX mult(IN1, IN2, design_res);
    assign design_is_correct = ((spec_res == design_res) ? 1 : 0);
    
endmodule



module WT_USP_RP_2x2_noX(
        input logic [1:0] IN1,
        input logic [1:0] IN2,
        output logic [3:0] result);
    
    
// Creating Partial Products 

    wire logic [1:0] pp0;
    wire logic [1:0] pp1;
    assign pp0 = {2{IN1[0]}} & IN2;
    assign pp1 = {2{IN1[1]}} & IN2;
    
    // The values to be summed in the summation tree, from LSB (left) to MSB:
     // pp0[0] pp0[1]   --   
     //   --   pp1[0] pp1[1] 
    
// Creating Summation Tree 

    
    assign result[0] = pp0[0];
    logic [2:0] adder_result;
    RP_2 final_adder ({pp1[1], pp0[1] }, {1'b0, pp1[0] }, adder_result );
    assign result[3:1] = adder_result[2:0];
endmodule



module RP_2 ( 
        input logic [1:0] IN1,
        input logic [1:0] IN2,
        output logic [2:0] OUT);
    
    logic C0, C1, C2;
    ha m0 (IN1[0], IN2[0], OUT[0], C0);
    fa m1 (IN1[1], IN2[1], C0, OUT[1], C1);
    assign OUT[2] = C1;

endmodule

module RP_2_spec (
        input logic [1:0] IN1,
        input logic [1:0] IN2,
        output logic adder_correct,
        output logic [2:0] spec_res);
    
    assign spec_res = IN1 + IN2;
    wire [2:0] adder_res;
    RP_2 adder(IN1, IN2, adder_res);
    assign adder_correct = ((spec_res == adder_res) ? 1 : 0);
    
endmodule



module ha (
        input logic a,
        input logic b,
        output logic s,
        output logic c);
    
    assign s = a ^ b;
    assign c = a & b;
endmodule



module fa (
        input logic x,
        input logic y,
        input logic z,
        output logic s,
        output logic c);
    
    assign s = x ^ y ^ z;
    assign c = (x & y) | (x & z) | (y & z);
endmodule

module Four2Two 
        #(parameter WIDTH=1) (
        input logic [WIDTH-1:0] in1,
        input logic [WIDTH-1:0] in2,
        input logic [WIDTH-1:0] in3,
        input logic [WIDTH-1:0] in4,
        input logic cin,
        output logic [WIDTH-1:0] sum,
        output logic [WIDTH-1:0] carry,
        output logic cout);
    
    wire logic [WIDTH:0] temp1;
    assign temp1 = {((in1 ^ in2)&in3 | in1 & ~(in1^in2)),cin};
    assign sum = ((in1 ^ in2) ^ in3 ^ in4) ^ temp1[WIDTH-1:0];
    assign carry = ((in1 ^ in2) ^ in3 ^ in4) & temp1[WIDTH-1:0] | in4 & ~((in1 ^ in2) ^ in3 ^ in4);
    assign cout = temp1[WIDTH];
endmodule




